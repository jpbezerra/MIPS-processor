cpu.dm.memory[0] = 8'b00000000;
cpu.dm.memory[1] = 8'b00000000;
cpu.dm.memory[2] = 8'b00000000;
cpu.dm.memory[3] = 8'b00000001;

cpu.dm.memory[4] = 8'b00000000;
cpu.dm.memory[5] = 8'b00000000;
cpu.dm.memory[6] = 8'b00000000;
cpu.dm.memory[7] = 8'b00000010;

cpu.dm.memory[8] = 8'b00000000;
cpu.dm.memory[9] = 8'b00000000;
cpu.dm.memory[10] = 8'b00000000;
cpu.dm.memory[11] = 8'b00000011;

cpu.dm.memory[12] = 8'b00000000;
cpu.dm.memory[13] = 8'b00000000;
cpu.dm.memory[14] = 8'b00000000;
cpu.dm.memory[15] = 8'b00000100;

cpu.dm.memory[16] = 8'b00000000;
cpu.dm.memory[17] = 8'b00000000;
cpu.dm.memory[18] = 8'b00000000;
cpu.dm.memory[19] = 8'b00000101;

cpu.dm.memory[20] = 8'b00000000;
cpu.dm.memory[21] = 8'b00000000;
cpu.dm.memory[22] = 8'b00000000;
cpu.dm.memory[23] = 8'b00000110;

cpu.dm.memory[24] = 8'b00000000;
cpu.dm.memory[25] = 8'b00000000;
cpu.dm.memory[26] = 8'b00000000;
cpu.dm.memory[27] = 8'b00000111;

cpu.dm.memory[28] = 8'b00000000;
cpu.dm.memory[29] = 8'b00000000;
cpu.dm.memory[30] = 8'b00000000;
cpu.dm.memory[31] = 8'b00001000;

